
module pool
(
    input max,
    input clk,
    input rst,
    input 
)

endmodule