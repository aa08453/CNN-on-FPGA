module tb_load_kernel();
    reg clk = 0;
    reg rst = 1;
    wire [7:0] k0, k1, k2, k3, k4, k5, k6, k7, k8;

    load_kernel uut (
        .clk(clk),
        .rst(rst),
        .kernel0(k0), .kernel1(k1), .kernel2(k2),
        .kernel3(k3), .kernel4(k4), .kernel5(k5),
        .kernel6(k6), .kernel7(k7), .kernel8(k8)
    );

    always #5 clk = ~clk;

    initial begin
        $dumpfile("w_load_kernel.vcd");
        $dumpvars(0, tb_load_kernel);

        #10 rst = 0;
        #20;

        $display("KERNEL:");
        $display("%d %d %d", k0, k1, k2);
        $display("%d %d %d", k3, k4, k5);
        $display("%d %d %d", k6, k7, k8);

        $finish;
    end
endmodule
